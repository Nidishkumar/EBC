// Module name: tb Module
// Module Description: Generating events for 16X16 pixel
// Author: [Your Name]
// Date: [Current Date]
// Version: [Version Number]
//------------------------------------------------------------------------------------------------------------------
import lib_arbiter_pkg::*;                                      // Importing arbiter package containing parameter constants

module tb_level;
  // Inputs
  logic clk_i                                   ; // Clock input
  logic reset_i                                 ; // Active high Reset input
  logic [ROWS-1:0][COLS-1:0][POLARITY-1:0]req_i;       // Request signals for each row and column, with POLARITY bits determining the signal's polarity or behavior
  // Outputs
 logic [ROWS-1:0][COLS-1:0] gnt_o             ; //grant output

 logic grp_release_o;
	logic [WIDTH-1:0] data_out_o;
  
  top_module
  dut (
            .clk_i        (clk_i)         ,     // Clock input
            .reset_i      (reset_i)       ,     // Active high Reset input
            .set_i        (req_i)         ,     // Request signals for each row and column, with POLARITY bits determining the signal's polarity 
            .gnt_o          (gnt_o)         ,     // grant outputs
				.grp_release_o(grp_release_o),
        .data_out_o(data_out_o)

  );


  // Clock generation
  initial begin
    clk_i = 0;
    forever #5 clk_i = ~clk_i; // Clock with a period of 10 time units
  end

  // Reset generation
  task apply_reset;
  begin
    reset_i = 1;
    #10 reset_i = 0;
  end
endtask
  //-------------------------------------------Deasserting request---------------------------------------------//

always_ff@(posedge clk_i)
 begin
 for(int i=0;i<ROWS;i++)
   begin
	 for(int j=0;j<ROWS;j++)
	  begin
	    if(gnt_o[i][j]==1'b1)
		   begin
		    req_i[i][j]<='0;
			end
	  end
	end 
end 
//----------------------------------------------Apply Request-------------------------------------------------------
task apply_request([ROWS-1:0][COLS-1:0][POLARITY-1:0]req);
begin
 req_i=req;
end
endtask
//-------------------------------------------End of Deasserting request---------------------------------------------//

  initial begin
    	 apply_reset;
	 //Random Events across pixel
   apply_request({
      {2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00}, // Row 0 inactive
      {2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01}, // Row 1 active
      {2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00}, // Row 2 inactive
      {2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b10, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10}, // Row 3 active
      {2'b01, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10}, // Row 4 inactive
      {2'b10, 2'b10, 2'b01, 2'b00, 2'b10, 2'b10, 2'b01, 2'b10, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b01}, // Row 5 active
      {2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00}, // Row 6 inactive
      {2'b01, 2'b01, 2'b10, 2'b10, 2'b10, 2'b01, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10}, // Row 7 active
      
		{2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00}, // Row 8 inactive
      {2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01}, // Row 9 active
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00}, // Row 10 inactive
      {2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b10}, // Row 11 active
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00}, // Row 12 inactive
      {2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b01}, // Row 13 active
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00}, // Row 14 inactive
      {2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10}  // Row 15 active
    });
	 #200;
	 
	 //  Alternate Row has Active events
	 apply_request({
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b10, 2'b10, 2'b01, 2'b00, 2'b10, 2'b10, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b00, 2'b10, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b10, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b10},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b01, 2'b01, 2'b01, 2'b10, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10, 2'b00, 2'b01, 2'b10, 2'b10, 2'b10, 2'b10},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b10, 2'b00},
		
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b01, 2'b01, 2'b01, 2'b10, 2'b10, 2'b10, 2'b01, 2'b01, 2'b01, 2'b10, 2'b00, 2'b01, 2'b01, 2'b10, 2'b10, 2'b10}
    });
	 #250;
	 apply_reset;
	  
	 //MSB 8rows of Pixel has active events
	  apply_request({
      {2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b00, 2'b10, 2'b00},
      {2'b00, 2'b10, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b10, 2'b00},
      {2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b10, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b10, 2'b01, 2'b10, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b01},
      {2'b10, 2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01},
      {2'b01, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b10, 2'b10, 2'b00, 2'b00, 2'b10},
      {2'b00, 2'b00, 2'b01, 2'b10, 2'b00, 2'b00, 2'b10, 2'b10, 2'b01, 2'b01, 2'b01, 2'b00, 2'b00, 2'b01, 2'b00, 2'b00},

      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
      {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
		{2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00}
		});
     
    #200;
	  //No activve Events 
	   apply_request( {
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00}
    });
	 
	 #200
	 //alternate pixel blocks has active events
	  apply_request({
        {2'b01, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b10, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b01, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00},
		  
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b10, 2'b10},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b10, 2'b10, 2'b01},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b10},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b01, 2'b10, 2'b01},
		  
        {2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b10, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b00, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
        {2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00},
		  
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b10, 2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b10, 2'b10, 2'b10},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b10, 2'b00, 2'b01},
        {2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b00, 2'b10}
    });
	 
	 #300;
	 //Active events 
	  apply_request({
	         {2'b10, 2'b10, 2'b01, 2'b00, 2'b00, 2'b01, 2'b10, 2'b10, 2'b10, 2'b01, 2'b01, 2'b10, 2'b01, 2'b00, 2'b10, 2'b00},
				{2'b01, 2'b00, 2'b10, 2'b10, 2'b10, 2'b01, 2'b10, 2'b01, 2'b01, 2'b00, 2'b10, 2'b10, 2'b00, 2'b10, 2'b10, 2'b01},
				{2'b10, 2'b00, 2'b00, 2'b00, 2'b00, 2'b10, 2'b00, 2'b00, 2'b10, 2'b01, 2'b01, 2'b00, 2'b10, 2'b01, 2'b01, 2'b10},
				{2'b01, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b01, 2'b01, 2'b01, 2'b10, 2'b10, 2'b10, 2'b01, 2'b10, 2'b00, 2'b10},
				
				{2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
				{2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
				{2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
				{2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
				
				{2'b01, 2'b00, 2'b01, 2'b00, 2'b01, 2'b10, 2'b00, 2'b10, 2'b10, 2'b01, 2'b01, 2'b01, 2'b01, 2'b01, 2'b00, 2'b10},
				{2'b10, 2'b10, 2'b00, 2'b01, 2'b10, 2'b00, 2'b01, 2'b00, 2'b10, 2'b10, 2'b00, 2'b10, 2'b00, 2'b10, 2'b01, 2'b00},
				{2'b01, 2'b10, 2'b10, 2'b10, 2'b10, 2'b00, 2'b10, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b00, 2'b10, 2'b10, 2'b00},
				{2'b01, 2'b01, 2'b01, 2'b00, 2'b01, 2'b10, 2'b10, 2'b00, 2'b01, 2'b01, 2'b00, 2'b01, 2'b01, 2'b01, 2'b10, 2'b10},
				
				{2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
				{2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
				{2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00},
				{2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00, 2'b00}
				});

	 $finish;
  end
endmodule