package arbiter_pkg;

  // Define parameters
  parameter ROWS = 8;
  parameter COLS = 8;
  parameter POLARITY = 2;
  parameter y_width = 3;
  parameter x_width = 3;
 
  parameter WIDTH = ROWS;
  parameter NUM_PORTS = WIDTH;


endpackage