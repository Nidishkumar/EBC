// Package:asyn_fifo_pkg
// Description: Centralized storage for parameters and constants used across design modules
// Date: 
// Version: 1.0
// Author: 

package asyn_fifo_pkg;

//synchronizer
//parameter int PTR_WIDTH = 3;

//wptr_handler
//parameter int PTR_WIDTH = 3;
//rptr_handler
//parameter int PTR_WIDTH = 3;
//fifo_mem 
parameter int DEPTH = 8;
parameter int DATA_WIDTH = 16;
parameter int PTR_WIDTH = 3;

//asynchronous_fifo
//parameter int DEPTH = 8;
//parameter int DATA_WIDTH = 8;
endpackage
