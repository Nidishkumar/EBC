// Module name: Polarity Selector Module
// Module Description: This Polarity Selector module outputs a selected polarity based on the request signals' polarity.
// Author: [Your Name]
// Date: [Current Date]
// Version: [Version Number]
//------------------------------------------------------------------------------------------------------------------

import lib_arbiter_pkg::*;  // Importing arbiter package containing parameter constants

// Define the module 'polarity_selector' with the following ports
module polarity_selector 
(
    input logic clk_i,              // Input clock signal (clk_i)
    input logic reset_i,            // Input reset signal (reset_i)
    input logic [POLARITY-1:0] req_i, // 2-bit input request signal (req_i)
    output logic polarity_out         // Output signal (polarity_out) representing the selected polarity
);

always_ff @(posedge clk_i or posedge reset_i) 
begin
    if (reset_i) 
    begin
        polarity_out <= 1'b0;  // Reset the output polarity to 0 when reset is triggered
    end
    else 
    begin
        // Case statement to determine the polarity output based on request signal (req_i)
        case(req_i)
            2'b10   : polarity_out <= 1'b1;  // If req_i is 2'b10, set polarity_out to 1,indicates intensity higher than threshold
            2'b01   : polarity_out <= 1'b0;  // If req_i is 2'b01, set polarity_out to 0,indicates intensity lower than threshold
            default : polarity_out <= 1'b0;  // Default case:set polarity_out to 0
        endcase
    end
end

endmodule



/*// Module name: Polarity Selecter Module
// Module Description: This Polarity Selecter module outputs based on polarity of requests.
// Author: [Your Name]
// Date: [Current Date]
// Version: [Version Number]
//------------------------------------------------------------------------------------------------------------------
import lib_arbiter_pkg::*;                   // Importing arbiter package containing parameter constants

module polarity_selector 

(
	input logic clk_i				  ,
	input logic reset_i				  ,
    input logic [POLARITY-1:0] req_i  ,     // 2-bit input request signal (req_i)
    output logic polarity_out               // Output signal (polarity_o) representing the selected polarity
);

 // Determine the polarity (pol_out) based on the request input (req_i) 

	always_ff @(posedge clk_i or posedge reset_i) 
	   begin
        if (reset_i) 
		   begin
				polarity_out <= 1'b0;
		   end
		else
	  		begin
				case(req_i)
					2'b10   :    polarity_out <= 1'b1;
					2'b01   :    polarity_out <= 1'b0;
					default :    polarity_out <= 1'b0;
				endcase
	  		end	 
	   end	 
endmodule */

  
  