// Package:syn_fifo_pkg
// Description: Centralized storage for parameters and constants used across design modules
// Date: 
// Version: 1.0
// Author: 

package syn_fifo_pkg;

parameter DEPTH=8;
parameter WIDTH=16;

endpackage
